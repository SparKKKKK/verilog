module fifo_ram(
wdata,rdata,waddr,raddr,write,read
    );