module fifo_ctrl(

    );